** Profile: "SCHEMATIC1-sim1"  [ D:\Ecole\EI-2I-3-S6\Electronique Analogique\TP\TP2\Pspce_TP2_julian_BARKOUDEH\tp2-schematic1-sim1.sim ] 

** Creating circuit file "tp2-schematic1-sim1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 50 10 100k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\tp2-SCHEMATIC1.net" 


.END
